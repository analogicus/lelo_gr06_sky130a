magic
tech sky130A
magscale 1 2
timestamp 1769081024
<< metal2 >>
rect 0 18989 400 19000
rect 0 18609 10 18989
rect 390 18609 400 18989
rect 0 890 400 18609
rect 0 510 10 890
rect 390 510 400 890
rect 0 0 400 510
rect 500 18490 900 19000
rect 500 18110 511 18490
rect 891 18110 900 18490
rect 500 390 900 18110
rect 500 10 510 390
rect 890 10 900 390
rect 500 0 900 10
rect 29100 18491 29500 19000
rect 29100 18111 29110 18491
rect 29490 18111 29500 18491
rect 29100 390 29500 18111
rect 29100 10 29110 390
rect 29490 10 29500 390
rect 29100 0 29500 10
rect 29600 18988 30000 19000
rect 29600 18608 29609 18988
rect 29989 18608 30000 18988
rect 29600 892 30000 18608
rect 29600 512 29611 892
rect 29991 512 30000 892
rect 29600 0 30000 512
<< via2 >>
rect 10 18609 390 18989
rect 10 510 390 890
rect 511 18110 891 18490
rect 510 10 890 390
rect 29110 18111 29490 18491
rect 29110 10 29490 390
rect 29609 18608 29989 18988
rect 29611 512 29991 892
<< metal3 >>
rect 0 18989 30000 19000
rect 0 18609 10 18989
rect 390 18988 30000 18989
rect 390 18609 29609 18988
rect 0 18608 29609 18609
rect 29989 18608 30000 18988
rect 0 18600 30000 18608
rect 0 18491 30000 18500
rect 0 18490 29110 18491
rect 0 18110 511 18490
rect 891 18111 29110 18490
rect 29490 18111 30000 18491
rect 891 18110 30000 18111
rect 0 18100 30000 18110
rect 6688 17618 6752 17624
rect 15528 17616 15534 17618
rect 6752 17556 15534 17616
rect 15528 17554 15534 17556
rect 15598 17554 15604 17618
rect 6688 17548 6752 17554
rect 0 892 30000 900
rect 0 890 29611 892
rect 0 510 10 890
rect 390 512 29611 890
rect 29991 512 30000 892
rect 390 510 30000 512
rect 0 500 30000 510
rect 0 390 30000 400
rect 0 10 510 390
rect 890 10 29110 390
rect 29490 10 30000 390
rect 0 0 30000 10
<< via3 >>
rect 6688 17554 6752 17618
rect 15534 17554 15598 17618
<< metal4 >>
rect 6690 18582 6750 19000
rect 6690 17619 6750 18502
rect 15522 18592 15582 19000
rect 15522 18413 15582 18512
rect 15522 18299 15596 18413
rect 15536 17619 15596 18299
rect 6687 17618 6753 17619
rect 6687 17554 6688 17618
rect 6752 17554 6753 17618
rect 6687 17553 6753 17554
rect 15533 17618 15599 17619
rect 15533 17554 15534 17618
rect 15598 17554 15599 17618
rect 15533 17553 15599 17554
<< rmetal4 >>
rect 6690 18502 6750 18582
rect 15522 18512 15582 18592
<< labels >>
flabel metal3 0 0 30000 400 0 FreeSans 1600 0 0 0 VSS
port 0 nsew signal input
flabel metal4 15522 18600 15582 19000 0 FreeSans 320 0 0 0 OSC_TEMP_1V8
port 1 nsew signal output
flabel metal4 6690 18599 6750 18999 0 FreeSans 320 0 0 0 PWRUP_1V8
port 2 nsew signal input
flabel metal3 0 18600 30000 19000 0 FreeSans 1600 0 0 0 VDD_1V8
port 3 nsew signal input
<< end >>
